`timescale 1ns / 1ps
// See LICENSE for licensing details.
module leopard_fpga
   (input wire aclk,
    input wire aresetn,
    input wire [7:0] ctrl_a,
    input wire [7:0] ctrl_i,
    output wire [7:0] ctrl_o);
    // instantiate Leopard root FPGA
endmodule: leopard_fpga